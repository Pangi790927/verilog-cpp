module mob();

endmodule