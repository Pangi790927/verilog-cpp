module cpu(
		A,
		B
	);
   
   input  A;
   output B;

   not(B, A);

endmodule